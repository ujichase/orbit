library ieee;
use ieee.std_logic_1164.all;

package const_pkg is

    constant FOO: std_logic := '0';

end package;