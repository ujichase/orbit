library ieee;
use ieee.std_logic_1164.all;

package a is

    constant MAGIC_KEY: std_logic_vector(31 downto 0) := x"CAFE_CAFE";

end package;