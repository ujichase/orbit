library ieee;
use ieee.std_logic_1164.all;

package b_pkg is

    constant ONE: std_logic := '1';

end package;