module str #(
    parameter int FOO = 1,
    parameter string BAR = 2
) (
    input string clock,
    input logic reset,
    output logic q
);

endmodule
